`ifndef INSTRUCTION_MEM
`define INSTRUCTION_MEM
`timescale 1ns / 1ps
module inst_mem(readaddr,instruction);
input [31:0]readaddr;
output [31:0] instruction;
reg [31:0]mem[127:0]; //size 128 words

//instruction load from where?

//initial begin
//$readmemb("C:/Users/Administrator/Desktop/VE370/Projects/project2/InstructionMem_for_P2_Demo.txt",mem);
//end
initial begin
//demo no bonus
mem[0]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[1]=32'b00100000000010010000000000110111 ;//addi $t1, $zero, 0x37
mem[2]=32'b00000001000010011000000000100100; //and $s0, $t0, $t1
mem[3]=32'b00000001000010011000000000100101; //or $s0, $t0, $t1
mem[4]=32'b10101100000100000000000000000100; //sw $s0, 4($zero)
mem[5]=32'b10101100000010000000000000001000; //sw $t0, 8($zero)
mem[6]=32'b00000001000010011000100000100000; //add $s1, $t0, $t1
mem[7]=32'b00000001000010011001000000100010; //sub $s2, $t0, $t1
mem[8]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[9]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[10]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[11]=32'b00010010001100100000000000010010; //beq $s1, $s2, error0
mem[12]=32'b10001100000100010000000000000100; //lw $s1, 4($zero)
mem[13]=32'b00110010001100100000000001001000; //andi $s2, $s1, 0x48
mem[14]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[15]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[16]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[17]=32'b00010010001100100000000000001111; //beq $s1, $s2, error1
mem[18]=32'b10001100000100110000000000001000; //lw $s3, 8($zero)
mem[19]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[20]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[21]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[22]=32'b00010010000100110000000000001101; //beq $s0, $s3, error2
mem[23]=32'b00000010010100011010000000101010; //slt $s4, $s2, $s1 (Last)
mem[24]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[25]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[26]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
mem[27]=32'b00010010100000000000000000001111; //beq $s4, $0, EXIT
mem[28]=32'b00000010001000001001000000100000; //add $s2, $s1, $0
mem[29]=32'b00001000000000000000000000010111; //j Last
mem[30]=32'b00100000000010000000000000000000;//addi $t0, $0, 0(error0)
mem[31]=32'b00100000000010010000000000000000; //addi $t1, $0, 0
mem[32]=32'b00001000000000000000000000111111; //j EXIT
mem[33]=32'b00100000000010000000000000000001; //addi $t0, $0, 1(error1)
mem[34]=32'b00100000000010010000000000000001; //addi $t1, $0, 1
mem[35]=32'b00001000000000000000000000111111; //j EXIT
mem[36]=32'b00100000000010000000000000000010; //addi $t0, $0, 2(error2)
mem[37]=32'b00100000000010010000000000000010; //addi $t1, $0, 2
mem[38]=32'b00001000000000000000000000111111; //j EXIT
mem[39]=32'b00100000000010000000000000000011; //addi $t0, $0, 3(error3)
mem[40]=32'b00100000000010010000000000000011; //addi $t1, $0, 3
mem[41]=32'b00001000000000000000000000111111; //j EXIT

//*************************
//bonus test
//mem[0]=32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
//mem[1]=32'b00100000000010010000000000110111 ;//addi $t1, $zero, 0x37
//mem[2]=32'b00000001000010011000000000100100; //and $s0, $t0, $t1
//mem[3]=32'b00000001000010011000000000100101; //or $s0, $t0, $t1
//mem[4]=32'b10101100000100000000000000000100; //sw $s0, 4($zero)
//mem[5]=32'b10101100000010000000000000001000; //sw $t0, 8($zero)
//mem[6]=32'b00000001000010011000100000100000; //add $s1, $t0, $t1
//mem[7]=32'b00000001000010011001000000100010; //sub $s2, $t0, $t1
//mem[8]=32'b00010010001100100000000000001001; //addi $t0, $zero, 0x20
//mem[9]=32'b10001100000100010000000000000100; //addi $t0, $zero, 0x20
//mem[10]=32'b00110010001100100000000001001000; //addi $t0, $zero, 0x20
//mem[11]=32'b00010010001100100000000000001001; //beq $s1, $s2, error0
//mem[12]=32'b10001100000100110000000000001000; //lw $s1, 4($zero)
//mem[13]=32'b00010010000100110000000000001010; //andi $s2, $s1, 0x48
//mem[14]=32'b00000010010100011010000000101010; //addi $t0, $zero, 0x20
//mem[15]=32'b00010010100000000000000000001111; //addi $t0, $zero, 0x20
//mem[16]=32'b00000010001000001001000000100000; //addi $t0, $zero, 0x20
//mem[17]=32'b00001000000000000000000000001110; //beq $s1, $s2, error1
//mem[18]=32'b00100000000010000000000000000000; //lw $s3, 8($zero)
//mem[19]=32'b00100000000010010000000000000000; //addi $t0, $zero, 0x20
//mem[20]=32'b00001000000000000000000000011111; //addi $t0, $zero, 0x20
//mem[21]=32'b00100000000010000000000000000001; //addi $t0, $zero, 0x20
//mem[22]=32'b00100000000010010000000000000001; //beq $s0, $s3, error2
//mem[23]=32'b00001000000000000000000000011111; //slt $s4, $s2, $s1 (Last)
//mem[24]=32'b00100000000010000000000000000010; //addi $t0, $zero, 0x20
//mem[25]=32'b00100000000010010000000000000010; //addi $t0, $zero, 0x20
//mem[26]=32'b00001000000000000000000000011111; //addi $t0, $zero, 0x20
//mem[27]=32'b00100000000010000000000000000011; //beq $s4, $0, EXIT
//mem[28]=32'b00100000000010010000000000000011; //add $s2, $s1, $0
//mem[29]=32'b00001000000000000000000000011111; //j Last


end
assign  instruction=mem[readaddr/4];


endmodule
`endif